magic
tech sky130A
magscale 1 2
timestamp 1745612919
<< viali >>
rect 4997 9129 5031 9163
rect 5365 9061 5399 9095
rect 1409 8993 1443 9027
rect 1685 8925 1719 8959
rect 2329 8925 2363 8959
rect 4813 8925 4847 8959
rect 5181 8925 5215 8959
rect 2513 8789 2547 8823
rect 1409 8449 1443 8483
rect 1593 8313 1627 8347
rect 4077 7905 4111 7939
rect 1409 7837 1443 7871
rect 1593 7837 1627 7871
rect 1869 7837 1903 7871
rect 3985 7837 4019 7871
rect 5181 7837 5215 7871
rect 1777 7701 1811 7735
rect 2053 7701 2087 7735
rect 4353 7701 4387 7735
rect 5365 7701 5399 7735
rect 4721 6953 4755 6987
rect 4813 6817 4847 6851
rect 1409 6749 1443 6783
rect 2697 6749 2731 6783
rect 4997 6749 5031 6783
rect 4721 6681 4755 6715
rect 1593 6613 1627 6647
rect 2881 6613 2915 6647
rect 5181 6613 5215 6647
rect 2789 6409 2823 6443
rect 5365 6409 5399 6443
rect 2973 6273 3007 6307
rect 4445 6273 4479 6307
rect 4721 6273 4755 6307
rect 5181 6273 5215 6307
rect 3157 6205 3191 6239
rect 4169 6205 4203 6239
rect 4537 6205 4571 6239
rect 3709 6137 3743 6171
rect 3801 6137 3835 6171
rect 4261 6137 4295 6171
rect 4445 6069 4479 6103
rect 4629 5865 4663 5899
rect 4537 5729 4571 5763
rect 4721 5661 4755 5695
rect 4813 5661 4847 5695
rect 1593 5321 1627 5355
rect 1409 5185 1443 5219
rect 5181 5185 5215 5219
rect 5365 4981 5399 5015
rect 4353 4777 4387 4811
rect 2329 4709 2363 4743
rect 4077 4641 4111 4675
rect 1501 4573 1535 4607
rect 2145 4573 2179 4607
rect 2513 4573 2547 4607
rect 2605 4573 2639 4607
rect 3985 4573 4019 4607
rect 4445 4573 4479 4607
rect 4629 4573 4663 4607
rect 1685 4437 1719 4471
rect 4537 4437 4571 4471
rect 3709 4233 3743 4267
rect 1409 4097 1443 4131
rect 2789 4097 2823 4131
rect 4077 4097 4111 4131
rect 5181 4097 5215 4131
rect 2881 4029 2915 4063
rect 3985 4029 4019 4063
rect 3157 3961 3191 3995
rect 1593 3893 1627 3927
rect 3893 3893 3927 3927
rect 5365 3893 5399 3927
rect 1869 3689 1903 3723
rect 1869 3485 1903 3519
rect 2053 3485 2087 3519
rect 1869 2601 1903 2635
rect 3801 2601 3835 2635
rect 1593 2533 1627 2567
rect 4077 2465 4111 2499
rect 4169 2465 4203 2499
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 3985 2397 4019 2431
rect 4261 2397 4295 2431
rect 4629 2397 4663 2431
rect 5089 2397 5123 2431
rect 5457 2329 5491 2363
rect 4813 2261 4847 2295
<< metal1 >>
rect 1104 9274 5796 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 5796 9274
rect 1104 9200 5796 9222
rect 4982 9120 4988 9172
rect 5040 9120 5046 9172
rect 5350 9052 5356 9104
rect 5408 9052 5414 9104
rect 1394 8984 1400 9036
rect 1452 8984 1458 9036
rect 1486 8916 1492 8968
rect 1544 8956 1550 8968
rect 1673 8959 1731 8965
rect 1673 8956 1685 8959
rect 1544 8928 1685 8956
rect 1544 8916 1550 8928
rect 1673 8925 1685 8928
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 2314 8916 2320 8968
rect 2372 8916 2378 8968
rect 4706 8916 4712 8968
rect 4764 8956 4770 8968
rect 4801 8959 4859 8965
rect 4801 8956 4813 8959
rect 4764 8928 4813 8956
rect 4764 8916 4770 8928
rect 4801 8925 4813 8928
rect 4847 8925 4859 8959
rect 4801 8919 4859 8925
rect 4890 8916 4896 8968
rect 4948 8956 4954 8968
rect 5169 8959 5227 8965
rect 5169 8956 5181 8959
rect 4948 8928 5181 8956
rect 4948 8916 4954 8928
rect 5169 8925 5181 8928
rect 5215 8925 5227 8959
rect 5169 8919 5227 8925
rect 1762 8780 1768 8832
rect 1820 8820 1826 8832
rect 2501 8823 2559 8829
rect 2501 8820 2513 8823
rect 1820 8792 2513 8820
rect 1820 8780 1826 8792
rect 2501 8789 2513 8792
rect 2547 8789 2559 8823
rect 2501 8783 2559 8789
rect 1104 8730 5796 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 5796 8730
rect 1104 8656 5796 8678
rect 842 8440 848 8492
rect 900 8480 906 8492
rect 1397 8483 1455 8489
rect 1397 8480 1409 8483
rect 900 8452 1409 8480
rect 900 8440 906 8452
rect 1397 8449 1409 8452
rect 1443 8449 1455 8483
rect 1397 8443 1455 8449
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 3878 8344 3884 8356
rect 1627 8316 3884 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 3878 8304 3884 8316
rect 3936 8304 3942 8356
rect 1104 8186 5796 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 5796 8186
rect 1104 8112 5796 8134
rect 4062 7896 4068 7948
rect 4120 7896 4126 7948
rect 1394 7828 1400 7880
rect 1452 7828 1458 7880
rect 1578 7828 1584 7880
rect 1636 7828 1642 7880
rect 1857 7871 1915 7877
rect 1857 7837 1869 7871
rect 1903 7837 1915 7871
rect 1857 7831 1915 7837
rect 1026 7760 1032 7812
rect 1084 7800 1090 7812
rect 1872 7800 1900 7831
rect 3970 7828 3976 7880
rect 4028 7828 4034 7880
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 5169 7871 5227 7877
rect 5169 7868 5181 7871
rect 4212 7840 5181 7868
rect 4212 7828 4218 7840
rect 5169 7837 5181 7840
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 1084 7772 1900 7800
rect 1084 7760 1090 7772
rect 1765 7735 1823 7741
rect 1765 7701 1777 7735
rect 1811 7732 1823 7735
rect 1854 7732 1860 7744
rect 1811 7704 1860 7732
rect 1811 7701 1823 7704
rect 1765 7695 1823 7701
rect 1854 7692 1860 7704
rect 1912 7692 1918 7744
rect 2041 7735 2099 7741
rect 2041 7701 2053 7735
rect 2087 7732 2099 7735
rect 4246 7732 4252 7744
rect 2087 7704 4252 7732
rect 2087 7701 2099 7704
rect 2041 7695 2099 7701
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 4341 7735 4399 7741
rect 4341 7701 4353 7735
rect 4387 7732 4399 7735
rect 5166 7732 5172 7744
rect 4387 7704 5172 7732
rect 4387 7701 4399 7704
rect 4341 7695 4399 7701
rect 5166 7692 5172 7704
rect 5224 7692 5230 7744
rect 5350 7692 5356 7744
rect 5408 7692 5414 7744
rect 1104 7642 5796 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 5796 7642
rect 1104 7568 5796 7590
rect 1104 7098 5796 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 5796 7098
rect 1104 7024 5796 7046
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 4709 6987 4767 6993
rect 4709 6984 4721 6987
rect 4304 6956 4721 6984
rect 4304 6944 4310 6956
rect 4709 6953 4721 6956
rect 4755 6953 4767 6987
rect 4709 6947 4767 6953
rect 3878 6808 3884 6860
rect 3936 6848 3942 6860
rect 4801 6851 4859 6857
rect 4801 6848 4813 6851
rect 3936 6820 4813 6848
rect 3936 6808 3942 6820
rect 4801 6817 4813 6820
rect 4847 6817 4859 6851
rect 4801 6811 4859 6817
rect 842 6740 848 6792
rect 900 6780 906 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 900 6752 1409 6780
rect 900 6740 906 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 2498 6740 2504 6792
rect 2556 6780 2562 6792
rect 2685 6783 2743 6789
rect 2685 6780 2697 6783
rect 2556 6752 2697 6780
rect 2556 6740 2562 6752
rect 2685 6749 2697 6752
rect 2731 6749 2743 6783
rect 4985 6783 5043 6789
rect 4985 6780 4997 6783
rect 2685 6743 2743 6749
rect 2792 6752 4997 6780
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 2406 6644 2412 6656
rect 1627 6616 2412 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 2406 6604 2412 6616
rect 2464 6644 2470 6656
rect 2792 6644 2820 6752
rect 4985 6749 4997 6752
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 3602 6672 3608 6724
rect 3660 6712 3666 6724
rect 4709 6715 4767 6721
rect 4709 6712 4721 6715
rect 3660 6684 4721 6712
rect 3660 6672 3666 6684
rect 4709 6681 4721 6684
rect 4755 6681 4767 6715
rect 4709 6675 4767 6681
rect 2464 6616 2820 6644
rect 2869 6647 2927 6653
rect 2464 6604 2470 6616
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 4154 6644 4160 6656
rect 2915 6616 4160 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 4614 6604 4620 6656
rect 4672 6644 4678 6656
rect 5169 6647 5227 6653
rect 5169 6644 5181 6647
rect 4672 6616 5181 6644
rect 4672 6604 4678 6616
rect 5169 6613 5181 6616
rect 5215 6613 5227 6647
rect 5169 6607 5227 6613
rect 1104 6554 5796 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 5796 6554
rect 1104 6480 5796 6502
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 2777 6443 2835 6449
rect 2777 6440 2789 6443
rect 2556 6412 2789 6440
rect 2556 6400 2562 6412
rect 2777 6409 2789 6412
rect 2823 6409 2835 6443
rect 2777 6403 2835 6409
rect 5350 6400 5356 6452
rect 5408 6400 5414 6452
rect 2958 6264 2964 6316
rect 3016 6264 3022 6316
rect 4430 6264 4436 6316
rect 4488 6264 4494 6316
rect 4614 6264 4620 6316
rect 4672 6304 4678 6316
rect 4709 6307 4767 6313
rect 4709 6304 4721 6307
rect 4672 6276 4721 6304
rect 4672 6264 4678 6276
rect 4709 6273 4721 6276
rect 4755 6273 4767 6307
rect 4709 6267 4767 6273
rect 4798 6264 4804 6316
rect 4856 6304 4862 6316
rect 5169 6307 5227 6313
rect 5169 6304 5181 6307
rect 4856 6276 5181 6304
rect 4856 6264 4862 6276
rect 5169 6273 5181 6276
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 3142 6196 3148 6248
rect 3200 6196 3206 6248
rect 4154 6196 4160 6248
rect 4212 6196 4218 6248
rect 4338 6196 4344 6248
rect 4396 6236 4402 6248
rect 4525 6239 4583 6245
rect 4525 6236 4537 6239
rect 4396 6208 4537 6236
rect 4396 6196 4402 6208
rect 4525 6205 4537 6208
rect 4571 6205 4583 6239
rect 4525 6199 4583 6205
rect 2314 6128 2320 6180
rect 2372 6168 2378 6180
rect 3697 6171 3755 6177
rect 3697 6168 3709 6171
rect 2372 6140 3709 6168
rect 2372 6128 2378 6140
rect 3697 6137 3709 6140
rect 3743 6137 3755 6171
rect 3697 6131 3755 6137
rect 3786 6128 3792 6180
rect 3844 6168 3850 6180
rect 4249 6171 4307 6177
rect 4249 6168 4261 6171
rect 3844 6140 4261 6168
rect 3844 6128 3850 6140
rect 4249 6137 4261 6140
rect 4295 6137 4307 6171
rect 4249 6131 4307 6137
rect 3050 6060 3056 6112
rect 3108 6100 3114 6112
rect 3970 6100 3976 6112
rect 3108 6072 3976 6100
rect 3108 6060 3114 6072
rect 3970 6060 3976 6072
rect 4028 6100 4034 6112
rect 4433 6103 4491 6109
rect 4433 6100 4445 6103
rect 4028 6072 4445 6100
rect 4028 6060 4034 6072
rect 4433 6069 4445 6072
rect 4479 6069 4491 6103
rect 4433 6063 4491 6069
rect 1104 6010 5796 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 5796 6010
rect 1104 5936 5796 5958
rect 2958 5856 2964 5908
rect 3016 5896 3022 5908
rect 4617 5899 4675 5905
rect 4617 5896 4629 5899
rect 3016 5868 4629 5896
rect 3016 5856 3022 5868
rect 4617 5865 4629 5868
rect 4663 5865 4675 5899
rect 4617 5859 4675 5865
rect 4246 5720 4252 5772
rect 4304 5760 4310 5772
rect 4522 5760 4528 5772
rect 4304 5732 4528 5760
rect 4304 5720 4310 5732
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 3602 5652 3608 5704
rect 3660 5692 3666 5704
rect 4709 5695 4767 5701
rect 4709 5692 4721 5695
rect 3660 5664 4721 5692
rect 3660 5652 3666 5664
rect 4709 5661 4721 5664
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5661 4859 5695
rect 4801 5655 4859 5661
rect 3878 5584 3884 5636
rect 3936 5624 3942 5636
rect 4816 5624 4844 5655
rect 3936 5596 4844 5624
rect 3936 5584 3942 5596
rect 1104 5466 5796 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 5796 5466
rect 1104 5392 5796 5414
rect 1394 5312 1400 5364
rect 1452 5352 1458 5364
rect 1581 5355 1639 5361
rect 1581 5352 1593 5355
rect 1452 5324 1593 5352
rect 1452 5312 1458 5324
rect 1581 5321 1593 5324
rect 1627 5352 1639 5355
rect 3970 5352 3976 5364
rect 1627 5324 3976 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 3970 5312 3976 5324
rect 4028 5352 4034 5364
rect 4430 5352 4436 5364
rect 4028 5324 4436 5352
rect 4028 5312 4034 5324
rect 4430 5312 4436 5324
rect 4488 5312 4494 5364
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 900 5188 1409 5216
rect 900 5176 906 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 4246 5176 4252 5228
rect 4304 5216 4310 5228
rect 5169 5219 5227 5225
rect 5169 5216 5181 5219
rect 4304 5188 5181 5216
rect 4304 5176 4310 5188
rect 5169 5185 5181 5188
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 1578 4972 1584 5024
rect 1636 5012 1642 5024
rect 4614 5012 4620 5024
rect 1636 4984 4620 5012
rect 1636 4972 1642 4984
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 5350 4972 5356 5024
rect 5408 4972 5414 5024
rect 1104 4922 5796 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 5796 4922
rect 1104 4848 5796 4870
rect 4341 4811 4399 4817
rect 4341 4777 4353 4811
rect 4387 4808 4399 4811
rect 4890 4808 4896 4820
rect 4387 4780 4896 4808
rect 4387 4777 4399 4780
rect 4341 4771 4399 4777
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 2317 4743 2375 4749
rect 2317 4709 2329 4743
rect 2363 4740 2375 4743
rect 4798 4740 4804 4752
rect 2363 4712 4804 4740
rect 2363 4709 2375 4712
rect 2317 4703 2375 4709
rect 4798 4700 4804 4712
rect 4856 4700 4862 4752
rect 3602 4672 3608 4684
rect 1504 4644 3608 4672
rect 1504 4616 1532 4644
rect 3602 4632 3608 4644
rect 3660 4672 3666 4684
rect 4065 4675 4123 4681
rect 4065 4672 4077 4675
rect 3660 4644 4077 4672
rect 3660 4632 3666 4644
rect 4065 4641 4077 4644
rect 4111 4641 4123 4675
rect 4065 4635 4123 4641
rect 1486 4564 1492 4616
rect 1544 4564 1550 4616
rect 1578 4564 1584 4616
rect 1636 4604 1642 4616
rect 2133 4607 2191 4613
rect 2133 4604 2145 4607
rect 1636 4576 2145 4604
rect 1636 4564 1642 4576
rect 2133 4573 2145 4576
rect 2179 4573 2191 4607
rect 2133 4567 2191 4573
rect 2406 4564 2412 4616
rect 2464 4604 2470 4616
rect 2501 4607 2559 4613
rect 2501 4604 2513 4607
rect 2464 4576 2513 4604
rect 2464 4564 2470 4576
rect 2501 4573 2513 4576
rect 2547 4573 2559 4607
rect 2501 4567 2559 4573
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4604 2651 4607
rect 3142 4604 3148 4616
rect 2639 4576 3148 4604
rect 2639 4573 2651 4576
rect 2593 4567 2651 4573
rect 3142 4564 3148 4576
rect 3200 4604 3206 4616
rect 3694 4604 3700 4616
rect 3200 4576 3700 4604
rect 3200 4564 3206 4576
rect 3694 4564 3700 4576
rect 3752 4564 3758 4616
rect 3878 4564 3884 4616
rect 3936 4604 3942 4616
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3936 4576 3985 4604
rect 3936 4564 3942 4576
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4430 4564 4436 4616
rect 4488 4564 4494 4616
rect 4614 4564 4620 4616
rect 4672 4564 4678 4616
rect 4706 4536 4712 4548
rect 1688 4508 4712 4536
rect 1688 4477 1716 4508
rect 4706 4496 4712 4508
rect 4764 4496 4770 4548
rect 1673 4471 1731 4477
rect 1673 4437 1685 4471
rect 1719 4437 1731 4471
rect 1673 4431 1731 4437
rect 4062 4428 4068 4480
rect 4120 4468 4126 4480
rect 4525 4471 4583 4477
rect 4525 4468 4537 4471
rect 4120 4440 4537 4468
rect 4120 4428 4126 4440
rect 4525 4437 4537 4440
rect 4571 4437 4583 4471
rect 4525 4431 4583 4437
rect 1104 4378 5796 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 5796 4378
rect 1104 4304 5796 4326
rect 3694 4224 3700 4276
rect 3752 4224 3758 4276
rect 842 4088 848 4140
rect 900 4128 906 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 900 4100 1409 4128
rect 900 4088 906 4100
rect 1397 4097 1409 4100
rect 1443 4097 1455 4131
rect 1397 4091 1455 4097
rect 2777 4131 2835 4137
rect 2777 4097 2789 4131
rect 2823 4128 2835 4131
rect 2958 4128 2964 4140
rect 2823 4100 2964 4128
rect 2823 4097 2835 4100
rect 2777 4091 2835 4097
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 3602 4088 3608 4140
rect 3660 4128 3666 4140
rect 4065 4131 4123 4137
rect 4065 4128 4077 4131
rect 3660 4100 4077 4128
rect 3660 4088 3666 4100
rect 4065 4097 4077 4100
rect 4111 4097 4123 4131
rect 4065 4091 4123 4097
rect 5166 4088 5172 4140
rect 5224 4088 5230 4140
rect 2869 4063 2927 4069
rect 2869 4029 2881 4063
rect 2915 4060 2927 4063
rect 3786 4060 3792 4072
rect 2915 4032 3792 4060
rect 2915 4029 2927 4032
rect 2869 4023 2927 4029
rect 3786 4020 3792 4032
rect 3844 4020 3850 4072
rect 3973 4063 4031 4069
rect 3973 4029 3985 4063
rect 4019 4060 4031 4063
rect 4522 4060 4528 4072
rect 4019 4032 4528 4060
rect 4019 4029 4031 4032
rect 3973 4023 4031 4029
rect 4522 4020 4528 4032
rect 4580 4020 4586 4072
rect 3145 3995 3203 4001
rect 3145 3961 3157 3995
rect 3191 3992 3203 3995
rect 5074 3992 5080 4004
rect 3191 3964 5080 3992
rect 3191 3961 3203 3964
rect 3145 3955 3203 3961
rect 5074 3952 5080 3964
rect 5132 3952 5138 4004
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 3050 3924 3056 3936
rect 1627 3896 3056 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 3050 3884 3056 3896
rect 3108 3884 3114 3936
rect 3878 3884 3884 3936
rect 3936 3884 3942 3936
rect 5350 3884 5356 3936
rect 5408 3884 5414 3936
rect 1104 3834 5796 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 5796 3834
rect 1104 3760 5796 3782
rect 1857 3723 1915 3729
rect 1857 3689 1869 3723
rect 1903 3720 1915 3723
rect 4246 3720 4252 3732
rect 1903 3692 4252 3720
rect 1903 3689 1915 3692
rect 1857 3683 1915 3689
rect 4246 3680 4252 3692
rect 4304 3680 4310 3732
rect 1854 3476 1860 3528
rect 1912 3476 1918 3528
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3516 2099 3519
rect 4062 3516 4068 3528
rect 2087 3488 4068 3516
rect 2087 3485 2099 3488
rect 2041 3479 2099 3485
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 1104 3290 5796 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 5796 3290
rect 1104 3216 5796 3238
rect 1104 2746 5796 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 5796 2746
rect 1104 2672 5796 2694
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 2958 2632 2964 2644
rect 1903 2604 2964 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 2958 2592 2964 2604
rect 3016 2592 3022 2644
rect 3789 2635 3847 2641
rect 3789 2601 3801 2635
rect 3835 2632 3847 2635
rect 4154 2632 4160 2644
rect 3835 2604 4160 2632
rect 3835 2601 3847 2604
rect 3789 2595 3847 2601
rect 4154 2592 4160 2604
rect 4212 2592 4218 2644
rect 4246 2592 4252 2644
rect 4304 2632 4310 2644
rect 4614 2632 4620 2644
rect 4304 2604 4620 2632
rect 4304 2592 4310 2604
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 1581 2567 1639 2573
rect 1581 2533 1593 2567
rect 1627 2564 1639 2567
rect 1627 2536 4292 2564
rect 1627 2533 1639 2536
rect 1581 2527 1639 2533
rect 3050 2456 3056 2508
rect 3108 2496 3114 2508
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3108 2468 4077 2496
rect 3108 2456 3114 2468
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 4065 2459 4123 2465
rect 4154 2456 4160 2508
rect 4212 2456 4218 2508
rect 842 2388 848 2440
rect 900 2428 906 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 900 2400 1409 2428
rect 900 2388 906 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 3970 2388 3976 2440
rect 4028 2388 4034 2440
rect 4264 2437 4292 2536
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2428 4307 2431
rect 4338 2428 4344 2440
rect 4295 2400 4344 2428
rect 4295 2397 4307 2400
rect 4249 2391 4307 2397
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 4617 2431 4675 2437
rect 4617 2397 4629 2431
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 1762 2320 1768 2372
rect 1820 2360 1826 2372
rect 4632 2360 4660 2391
rect 5074 2388 5080 2440
rect 5132 2388 5138 2440
rect 1820 2332 4660 2360
rect 1820 2320 1826 2332
rect 5442 2320 5448 2372
rect 5500 2320 5506 2372
rect 4798 2252 4804 2304
rect 4856 2252 4862 2304
rect 1104 2202 5796 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 5796 2202
rect 1104 2128 5796 2150
<< via1 >>
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 4988 9163 5040 9172
rect 4988 9129 4997 9163
rect 4997 9129 5031 9163
rect 5031 9129 5040 9163
rect 4988 9120 5040 9129
rect 5356 9095 5408 9104
rect 5356 9061 5365 9095
rect 5365 9061 5399 9095
rect 5399 9061 5408 9095
rect 5356 9052 5408 9061
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 1492 8916 1544 8968
rect 2320 8959 2372 8968
rect 2320 8925 2329 8959
rect 2329 8925 2363 8959
rect 2363 8925 2372 8959
rect 2320 8916 2372 8925
rect 4712 8916 4764 8968
rect 4896 8916 4948 8968
rect 1768 8780 1820 8832
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 848 8440 900 8492
rect 3884 8304 3936 8356
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 4068 7939 4120 7948
rect 4068 7905 4077 7939
rect 4077 7905 4111 7939
rect 4111 7905 4120 7939
rect 4068 7896 4120 7905
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 1032 7760 1084 7812
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 4160 7828 4212 7880
rect 1860 7692 1912 7744
rect 4252 7692 4304 7744
rect 5172 7692 5224 7744
rect 5356 7735 5408 7744
rect 5356 7701 5365 7735
rect 5365 7701 5399 7735
rect 5399 7701 5408 7735
rect 5356 7692 5408 7701
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 4252 6944 4304 6996
rect 3884 6808 3936 6860
rect 848 6740 900 6792
rect 2504 6740 2556 6792
rect 2412 6604 2464 6656
rect 3608 6672 3660 6724
rect 4160 6604 4212 6656
rect 4620 6604 4672 6656
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 2504 6400 2556 6452
rect 5356 6443 5408 6452
rect 5356 6409 5365 6443
rect 5365 6409 5399 6443
rect 5399 6409 5408 6443
rect 5356 6400 5408 6409
rect 2964 6307 3016 6316
rect 2964 6273 2973 6307
rect 2973 6273 3007 6307
rect 3007 6273 3016 6307
rect 2964 6264 3016 6273
rect 4436 6307 4488 6316
rect 4436 6273 4445 6307
rect 4445 6273 4479 6307
rect 4479 6273 4488 6307
rect 4436 6264 4488 6273
rect 4620 6264 4672 6316
rect 4804 6264 4856 6316
rect 3148 6239 3200 6248
rect 3148 6205 3157 6239
rect 3157 6205 3191 6239
rect 3191 6205 3200 6239
rect 3148 6196 3200 6205
rect 4160 6239 4212 6248
rect 4160 6205 4169 6239
rect 4169 6205 4203 6239
rect 4203 6205 4212 6239
rect 4160 6196 4212 6205
rect 4344 6196 4396 6248
rect 2320 6128 2372 6180
rect 3792 6171 3844 6180
rect 3792 6137 3801 6171
rect 3801 6137 3835 6171
rect 3835 6137 3844 6171
rect 3792 6128 3844 6137
rect 3056 6060 3108 6112
rect 3976 6060 4028 6112
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 2964 5856 3016 5908
rect 4252 5720 4304 5772
rect 4528 5763 4580 5772
rect 4528 5729 4537 5763
rect 4537 5729 4571 5763
rect 4571 5729 4580 5763
rect 4528 5720 4580 5729
rect 3608 5652 3660 5704
rect 3884 5584 3936 5636
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 1400 5312 1452 5364
rect 3976 5312 4028 5364
rect 4436 5312 4488 5364
rect 848 5176 900 5228
rect 4252 5176 4304 5228
rect 1584 4972 1636 5024
rect 4620 4972 4672 5024
rect 5356 5015 5408 5024
rect 5356 4981 5365 5015
rect 5365 4981 5399 5015
rect 5399 4981 5408 5015
rect 5356 4972 5408 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 4896 4768 4948 4820
rect 4804 4700 4856 4752
rect 3608 4632 3660 4684
rect 1492 4607 1544 4616
rect 1492 4573 1501 4607
rect 1501 4573 1535 4607
rect 1535 4573 1544 4607
rect 1492 4564 1544 4573
rect 1584 4564 1636 4616
rect 2412 4564 2464 4616
rect 3148 4564 3200 4616
rect 3700 4564 3752 4616
rect 3884 4564 3936 4616
rect 4436 4607 4488 4616
rect 4436 4573 4445 4607
rect 4445 4573 4479 4607
rect 4479 4573 4488 4607
rect 4436 4564 4488 4573
rect 4620 4607 4672 4616
rect 4620 4573 4629 4607
rect 4629 4573 4663 4607
rect 4663 4573 4672 4607
rect 4620 4564 4672 4573
rect 4712 4496 4764 4548
rect 4068 4428 4120 4480
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 3700 4267 3752 4276
rect 3700 4233 3709 4267
rect 3709 4233 3743 4267
rect 3743 4233 3752 4267
rect 3700 4224 3752 4233
rect 848 4088 900 4140
rect 2964 4088 3016 4140
rect 3608 4088 3660 4140
rect 5172 4131 5224 4140
rect 5172 4097 5181 4131
rect 5181 4097 5215 4131
rect 5215 4097 5224 4131
rect 5172 4088 5224 4097
rect 3792 4020 3844 4072
rect 4528 4020 4580 4072
rect 5080 3952 5132 4004
rect 3056 3884 3108 3936
rect 3884 3927 3936 3936
rect 3884 3893 3893 3927
rect 3893 3893 3927 3927
rect 3927 3893 3936 3927
rect 3884 3884 3936 3893
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 4252 3680 4304 3732
rect 1860 3519 1912 3528
rect 1860 3485 1869 3519
rect 1869 3485 1903 3519
rect 1903 3485 1912 3519
rect 1860 3476 1912 3485
rect 4068 3476 4120 3528
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 2964 2592 3016 2644
rect 4160 2592 4212 2644
rect 4252 2592 4304 2644
rect 4620 2592 4672 2644
rect 3056 2456 3108 2508
rect 4160 2499 4212 2508
rect 4160 2465 4169 2499
rect 4169 2465 4203 2499
rect 4203 2465 4212 2499
rect 4160 2456 4212 2465
rect 848 2388 900 2440
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 3976 2431 4028 2440
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 4344 2388 4396 2440
rect 1768 2320 1820 2372
rect 5080 2431 5132 2440
rect 5080 2397 5089 2431
rect 5089 2397 5123 2431
rect 5123 2397 5132 2431
rect 5080 2388 5132 2397
rect 5448 2363 5500 2372
rect 5448 2329 5457 2363
rect 5457 2329 5491 2363
rect 5491 2329 5500 2363
rect 5448 2320 5500 2329
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
<< metal2 >>
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 4986 10432 5042 10441
rect 4986 10367 5042 10376
rect 1412 9042 1440 10367
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 5000 9178 5028 10367
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5356 9104 5408 9110
rect 5354 9072 5356 9081
rect 5408 9072 5410 9081
rect 1400 9036 1452 9042
rect 5354 9007 5410 9016
rect 1400 8978 1452 8984
rect 1492 8968 1544 8974
rect 846 8936 902 8945
rect 1492 8910 1544 8916
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 846 8871 902 8880
rect 860 8498 888 8871
rect 848 8492 900 8498
rect 848 8434 900 8440
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1032 7812 1084 7818
rect 1032 7754 1084 7760
rect 1044 7721 1072 7754
rect 1030 7712 1086 7721
rect 1030 7647 1086 7656
rect 848 6792 900 6798
rect 848 6734 900 6740
rect 860 6497 888 6734
rect 846 6488 902 6497
rect 846 6423 902 6432
rect 1412 5370 1440 7822
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 860 5137 888 5170
rect 846 5128 902 5137
rect 846 5063 902 5072
rect 1504 4622 1532 8910
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1596 5030 1624 7822
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1596 4622 1624 4966
rect 1492 4616 1544 4622
rect 1492 4558 1544 4564
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 848 4140 900 4146
rect 848 4082 900 4088
rect 860 3777 888 4082
rect 846 3768 902 3777
rect 846 3703 902 3712
rect 848 2440 900 2446
rect 846 2408 848 2417
rect 1676 2440 1728 2446
rect 900 2408 902 2417
rect 1676 2382 1728 2388
rect 846 2343 902 2352
rect 1688 921 1716 2382
rect 1780 2378 1808 8774
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1872 3534 1900 7686
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 2332 6186 2360 8910
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 3884 8356 3936 8362
rect 3884 8298 3936 8304
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 3896 6866 3924 8298
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2320 6180 2372 6186
rect 2320 6122 2372 6128
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2424 4622 2452 6598
rect 2516 6458 2544 6734
rect 3608 6724 3660 6730
rect 3608 6666 3660 6672
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2976 5914 3004 6258
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2976 2650 3004 4082
rect 3068 3942 3096 6054
rect 3160 4622 3188 6190
rect 3620 5710 3648 6666
rect 3792 6180 3844 6186
rect 3792 6122 3844 6128
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 3620 4690 3648 5646
rect 3608 4684 3660 4690
rect 3608 4626 3660 4632
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3620 4146 3648 4626
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3712 4282 3740 4558
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3804 4078 3832 6122
rect 3896 5642 3924 6802
rect 3988 6118 4016 7822
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 3896 4622 3924 5578
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3896 3942 3924 4558
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3068 2514 3096 3878
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 3988 2446 4016 5306
rect 4080 4486 4108 7890
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4172 6662 4200 7822
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4264 7002 4292 7686
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 4080 3534 4108 4422
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4172 2650 4200 6190
rect 4264 5778 4292 6938
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4632 6322 4660 6598
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 4264 3738 4292 5170
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4264 2530 4292 2586
rect 4172 2514 4292 2530
rect 4160 2508 4292 2514
rect 4212 2502 4292 2508
rect 4160 2450 4212 2456
rect 4356 2446 4384 6190
rect 4448 5370 4476 6258
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4448 4622 4476 5306
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 4540 4078 4568 5714
rect 4632 5030 4660 6258
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4632 4622 4660 4966
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4632 2650 4660 4558
rect 4724 4554 4752 8910
rect 4804 6316 4856 6322
rect 4804 6258 4856 6264
rect 4816 4758 4844 6258
rect 4908 4826 4936 8910
rect 5172 7744 5224 7750
rect 5356 7744 5408 7750
rect 5172 7686 5224 7692
rect 5354 7712 5356 7721
rect 5408 7712 5410 7721
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 5184 4146 5212 7686
rect 5354 7647 5410 7656
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5368 6361 5396 6394
rect 5354 6352 5410 6361
rect 5354 6287 5410 6296
rect 5356 5024 5408 5030
rect 5354 4992 5356 5001
rect 5408 4992 5410 5001
rect 5354 4927 5410 4936
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5080 4004 5132 4010
rect 5080 3946 5132 3952
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 5092 2446 5120 3946
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5368 3641 5396 3878
rect 5354 3632 5410 3641
rect 5354 3567 5410 3576
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 5080 2440 5132 2446
rect 5080 2382 5132 2388
rect 1768 2372 1820 2378
rect 1768 2314 1820 2320
rect 5448 2372 5500 2378
rect 5448 2314 5500 2320
rect 4804 2304 4856 2310
rect 4802 2272 4804 2281
rect 4856 2272 4858 2281
rect 2610 2204 2918 2213
rect 4802 2207 4858 2216
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 5460 921 5488 2314
rect 1674 912 1730 921
rect 1674 847 1730 856
rect 5446 912 5502 921
rect 5446 847 5502 856
<< via2 >>
rect 1398 10376 1454 10432
rect 4986 10376 5042 10432
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 5354 9052 5356 9072
rect 5356 9052 5408 9072
rect 5408 9052 5410 9072
rect 5354 9016 5410 9052
rect 846 8880 902 8936
rect 1030 7656 1086 7712
rect 846 6432 902 6488
rect 846 5072 902 5128
rect 846 3712 902 3768
rect 846 2388 848 2408
rect 848 2388 900 2408
rect 900 2388 902 2408
rect 846 2352 902 2388
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 5354 7692 5356 7712
rect 5356 7692 5408 7712
rect 5408 7692 5410 7712
rect 5354 7656 5410 7692
rect 5354 6296 5410 6352
rect 5354 4972 5356 4992
rect 5356 4972 5408 4992
rect 5408 4972 5410 4992
rect 5354 4936 5410 4972
rect 5354 3576 5410 3632
rect 4802 2252 4804 2272
rect 4804 2252 4856 2272
rect 4856 2252 4858 2272
rect 4802 2216 4858 2252
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 1674 856 1730 912
rect 5446 856 5502 912
<< metal3 >>
rect 0 10434 800 10464
rect 1393 10434 1459 10437
rect 0 10432 1459 10434
rect 0 10376 1398 10432
rect 1454 10376 1459 10432
rect 0 10374 1459 10376
rect 0 10344 800 10374
rect 1393 10371 1459 10374
rect 4981 10434 5047 10437
rect 6100 10434 6900 10464
rect 4981 10432 6900 10434
rect 4981 10376 4986 10432
rect 5042 10376 6900 10432
rect 4981 10374 6900 10376
rect 4981 10371 5047 10374
rect 6100 10344 6900 10374
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 0 9074 800 9104
rect 5349 9074 5415 9077
rect 6100 9074 6900 9104
rect 0 8984 858 9074
rect 5349 9072 6900 9074
rect 5349 9016 5354 9072
rect 5410 9016 6900 9072
rect 5349 9014 6900 9016
rect 5349 9011 5415 9014
rect 6100 8984 6900 9014
rect 798 8941 858 8984
rect 798 8936 907 8941
rect 798 8880 846 8936
rect 902 8880 907 8936
rect 798 8878 907 8880
rect 841 8875 907 8878
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 0 7714 800 7744
rect 1025 7714 1091 7717
rect 0 7712 1091 7714
rect 0 7656 1030 7712
rect 1086 7656 1091 7712
rect 0 7654 1091 7656
rect 0 7624 800 7654
rect 1025 7651 1091 7654
rect 5349 7714 5415 7717
rect 6100 7714 6900 7744
rect 5349 7712 6900 7714
rect 5349 7656 5354 7712
rect 5410 7656 6900 7712
rect 5349 7654 6900 7656
rect 5349 7651 5415 7654
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 6100 7624 6900 7654
rect 2606 7583 2922 7584
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 841 6490 907 6493
rect 798 6488 907 6490
rect 798 6432 846 6488
rect 902 6432 907 6488
rect 798 6427 907 6432
rect 798 6384 858 6427
rect 0 6294 858 6384
rect 5349 6354 5415 6357
rect 6100 6354 6900 6384
rect 5349 6352 6900 6354
rect 5349 6296 5354 6352
rect 5410 6296 6900 6352
rect 5349 6294 6900 6296
rect 0 6264 800 6294
rect 5349 6291 5415 6294
rect 6100 6264 6900 6294
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 841 5130 907 5133
rect 798 5128 907 5130
rect 798 5072 846 5128
rect 902 5072 907 5128
rect 798 5067 907 5072
rect 798 5024 858 5067
rect 0 4934 858 5024
rect 5349 4994 5415 4997
rect 6100 4994 6900 5024
rect 5349 4992 6900 4994
rect 5349 4936 5354 4992
rect 5410 4936 6900 4992
rect 5349 4934 6900 4936
rect 0 4904 800 4934
rect 5349 4931 5415 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 6100 4904 6900 4934
rect 1946 4863 2262 4864
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 841 3770 907 3773
rect 798 3768 907 3770
rect 798 3712 846 3768
rect 902 3712 907 3768
rect 798 3707 907 3712
rect 798 3664 858 3707
rect 0 3574 858 3664
rect 5349 3634 5415 3637
rect 6100 3634 6900 3664
rect 5349 3632 6900 3634
rect 5349 3576 5354 3632
rect 5410 3576 6900 3632
rect 5349 3574 6900 3576
rect 0 3544 800 3574
rect 5349 3571 5415 3574
rect 6100 3544 6900 3574
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 841 2410 907 2413
rect 798 2408 907 2410
rect 798 2352 846 2408
rect 902 2352 907 2408
rect 798 2347 907 2352
rect 798 2304 858 2347
rect 0 2214 858 2304
rect 4797 2274 4863 2277
rect 6100 2274 6900 2304
rect 4797 2272 6900 2274
rect 4797 2216 4802 2272
rect 4858 2216 6900 2272
rect 4797 2214 6900 2216
rect 0 2184 800 2214
rect 4797 2211 4863 2214
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 6100 2184 6900 2214
rect 2606 2143 2922 2144
rect 0 914 800 944
rect 1669 914 1735 917
rect 0 912 1735 914
rect 0 856 1674 912
rect 1730 856 1735 912
rect 0 854 1735 856
rect 0 824 800 854
rect 1669 851 1735 854
rect 5441 914 5507 917
rect 6100 914 6900 944
rect 5441 912 6900 914
rect 5441 856 5446 912
rect 5502 856 6900 912
rect 5441 854 6900 856
rect 5441 851 5507 854
rect 6100 824 6900 854
<< via3 >>
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
<< metal4 >>
rect 1944 9280 2264 9296
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8192 2264 9216
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 8736 2924 9296
rect 2604 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3296 2924 4320
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
use sky130_fd_sc_hd__or4_2  _09_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4692 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _10_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _11_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _12_
timestamp 1704896540
transform 1 0 1840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _13_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _14_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _15_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4784 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _16_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4232 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _17_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2576 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _18_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2576 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _19_
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _20_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4140 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _21_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _22_
timestamp 1704896540
transform -1 0 3220 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 1704896540
transform -1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _24_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 1704896540
transform -1 0 1748 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_36 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4416 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_39 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4692 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_47
timestamp 1704896540
transform 1 0 5428 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_7
timestamp 1704896540
transform 1 0 1748 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_11
timestamp 1704896540
transform 1 0 2116 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_23
timestamp 1704896540
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_47
timestamp 1704896540
transform 1 0 5428 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_6
timestamp 1704896540
transform 1 0 1656 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_14
timestamp 1704896540
transform 1 0 2392 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_23
timestamp 1704896540
transform 1 0 3220 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3588 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_33
timestamp 1704896540
transform 1 0 4140 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_7
timestamp 1704896540
transform 1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_17
timestamp 1704896540
transform 1 0 2668 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_25
timestamp 1704896540
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_39
timestamp 1704896540
transform 1 0 4692 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_47
timestamp 1704896540
transform 1 0 5428 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_6
timestamp 1704896540
transform 1 0 1656 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_18
timestamp 1704896540
transform 1 0 2760 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_30
timestamp 1704896540
transform 1 0 3864 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_42
timestamp 1704896540
transform 1 0 4968 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1704896540
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_47
timestamp 1704896540
transform 1 0 5428 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_15
timestamp 1704896540
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_23
timestamp 1704896540
transform 1 0 3220 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3588 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_40
timestamp 1704896540
transform 1 0 4784 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_6
timestamp 1704896540
transform 1 0 1656 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_14
timestamp 1704896540
transform 1 0 2392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_20
timestamp 1704896540
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_37
timestamp 1704896540
transform 1 0 4508 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_46
timestamp 1704896540
transform 1 0 5336 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1704896540
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1704896540
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_39
timestamp 1704896540
transform 1 0 4692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_47
timestamp 1704896540
transform 1 0 5428 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_11
timestamp 1704896540
transform 1 0 2116 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_23
timestamp 1704896540
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1704896540
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_36
timestamp 1704896540
transform 1 0 4416 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_6
timestamp 1704896540
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_18
timestamp 1704896540
transform 1 0 2760 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_30
timestamp 1704896540
transform 1 0 3864 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_42
timestamp 1704896540
transform 1 0 4968 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_16
timestamp 1704896540
transform 1 0 2576 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_37
timestamp 1704896540
transform 1 0 4508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1704896540
transform 1 0 1840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1704896540
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1704896540
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1704896540
transform -1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1704896540
transform 1 0 5152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1704896540
transform 1 0 5152 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1704896540
transform 1 0 5152 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1704896540
transform 1 0 5152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1704896540
transform 1 0 5152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1704896540
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_13
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_14
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_15
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_16
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_17
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_18
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_19
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 5796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_20
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_21
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 5796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_22
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_23
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 5796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_24
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_25
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_27
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_28
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_29
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_30
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_31
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_32
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
<< labels >>
flabel metal4 s 2604 2128 2924 9296 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1944 2128 2264 9296 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 in[0]
port 2 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 in[1]
port 3 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 in[2]
port 4 nsew signal input
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 in[3]
port 5 nsew signal input
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 in[4]
port 6 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 in[5]
port 7 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 in[6]
port 8 nsew signal input
flabel metal3 s 0 824 800 944 0 FreeSans 480 0 0 0 in[7]
port 9 nsew signal input
flabel metal3 s 6100 10344 6900 10464 0 FreeSans 480 0 0 0 out[0]
port 10 nsew signal output
flabel metal3 s 6100 8984 6900 9104 0 FreeSans 480 0 0 0 out[1]
port 11 nsew signal output
flabel metal3 s 6100 7624 6900 7744 0 FreeSans 480 0 0 0 out[2]
port 12 nsew signal output
flabel metal3 s 6100 6264 6900 6384 0 FreeSans 480 0 0 0 out[3]
port 13 nsew signal output
flabel metal3 s 6100 4904 6900 5024 0 FreeSans 480 0 0 0 out[4]
port 14 nsew signal output
flabel metal3 s 6100 3544 6900 3664 0 FreeSans 480 0 0 0 out[5]
port 15 nsew signal output
flabel metal3 s 6100 2184 6900 2304 0 FreeSans 480 0 0 0 out[6]
port 16 nsew signal output
flabel metal3 s 6100 824 6900 944 0 FreeSans 480 0 0 0 out[7]
port 17 nsew signal output
rlabel metal1 3450 8704 3450 8704 0 VGND
rlabel metal1 3450 9248 3450 9248 0 VPWR
rlabel metal1 1886 4590 1886 4590 0 _00_
rlabel metal1 4324 4454 4324 4454 0 _01_
rlabel metal1 1840 7718 1840 7718 0 _02_
rlabel metal1 4002 2618 4002 2618 0 _03_
rlabel metal2 3818 5100 3818 5100 0 _04_
rlabel metal1 3036 6154 3036 6154 0 _05_
rlabel via1 3174 4590 3174 4590 0 _06_
rlabel metal1 3818 5882 3818 5882 0 _07_
rlabel metal1 2668 6426 2668 6426 0 _08_
rlabel metal3 1050 10404 1050 10404 0 in[0]
rlabel metal3 751 9044 751 9044 0 in[1]
rlabel metal3 866 7684 866 7684 0 in[2]
rlabel metal3 751 6324 751 6324 0 in[3]
rlabel metal3 751 4964 751 4964 0 in[4]
rlabel metal3 751 3604 751 3604 0 in[5]
rlabel metal3 751 2244 751 2244 0 in[6]
rlabel metal3 1188 884 1188 884 0 in[7]
rlabel metal1 2806 4658 2806 4658 0 net1
rlabel metal1 4646 4794 4646 4794 0 net10
rlabel metal1 3542 6630 3542 6630 0 net11
rlabel metal1 3588 4726 3588 4726 0 net12
rlabel metal1 3082 3706 3082 3706 0 net13
rlabel metal1 4784 7718 4784 7718 0 net14
rlabel metal1 3220 2346 3220 2346 0 net15
rlabel metal2 5106 3196 5106 3196 0 net16
rlabel metal1 4370 6834 4370 6834 0 net2
rlabel metal2 4554 4896 4554 4896 0 net3
rlabel metal1 2208 6630 2208 6630 0 net4
rlabel metal1 1518 5338 1518 5338 0 net5
rlabel metal1 2346 3910 2346 3910 0 net6
rlabel metal1 4324 2414 4324 2414 0 net7
rlabel metal1 2438 2618 2438 2618 0 net8
rlabel metal1 1702 4488 1702 4488 0 net9
rlabel metal2 5014 9775 5014 9775 0 out[0]
rlabel via2 5382 9061 5382 9061 0 out[1]
rlabel via2 5382 7701 5382 7701 0 out[2]
rlabel metal2 5382 6375 5382 6375 0 out[3]
rlabel via2 5382 4981 5382 4981 0 out[4]
rlabel metal2 5382 3757 5382 3757 0 out[5]
rlabel via2 4830 2261 4830 2261 0 out[6]
rlabel metal2 5474 1615 5474 1615 0 out[7]
<< properties >>
string FIXED_BBOX 0 0 6900 11424
<< end >>
